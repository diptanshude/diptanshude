module rca_4bit_20BEE0016(
    input [3:0] a,b,
    input cin,
    output [4:0] s
    );
    
    wire [3:0] w ;
    fa_df fa1(a[0],b[0],cin,s[0],w[1]);
    fa_df fa2(a[1],b[1],w[1],s[1],w[2]);
    fa_df fa3(a[2],b[2],w[2],s[2],w[3]);
    fa_df fa4(a[3],b[3],w[3],s[3],s[4]);
    
endmodule
   
module fa_df(
    input a,b,cin,
    output s,cout
    );
    
   assign s = a^b^cin;
   assign cout = (a&b)|(b&cin)|(a&cin);
   
endmodule
